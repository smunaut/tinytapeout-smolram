/*
 * user_module_341426151397261906.v
 */

`default_nettype none

module user_module_341426151397261906 (
	input  wire  [7:0] io_in,
	output wire  [7:0] io_out
);

	assign io_out = io_in;

endmodule // user_module_341426151397261906
